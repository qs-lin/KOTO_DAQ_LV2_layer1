-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 9.1 Build 222 10/21/2009 SJ Full Version"
-- CREATED		"Wed Sep 16 11:31:28 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY word_aligner IS 
	PORT
	(
		reset :  IN  STD_LOGIC;
		enable :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		buffer_data :  IN  STD_LOGIC_VECTOR(223 DOWNTO 0);
		compr_mask :  IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		out :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END word_aligner;

ARCHITECTURE bdf_type OF word_aligner IS 

COMPONENT and16
	PORT(data0x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT or16b
	PORT(data : IN STD_LOGIC_VECTOR(15 DOWNTO 0 , 0 TO 0);
		 result : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT and4b
	PORT(data : IN STD_LOGIC_VECTOR(3 DOWNTO 0 , 0 TO 0);
		 result : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT and3b
	PORT(data : IN STD_LOGIC_VECTOR(2 DOWNTO 0 , 0 TO 0);
		 result : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT and2b
	PORT(data : IN STD_LOGIC_VECTOR(1 DOWNTO 0 , 0 TO 0);
		 result : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT or15b
	PORT(data : IN STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
		 result : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT inv16b
	PORT(data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT inv1
	PORT(data : IN STD_LOGIC;
		 result : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT reg13set
	PORT(sset : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 aset : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const2
	PORT(		 result : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT or8b
	PORT(data : IN STD_LOGIC_VECTOR(7 DOWNTO 0 , 0 TO 0);
		 result : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT or12b
	PORT(data : IN STD_LOGIC_VECTOR(11 DOWNTO 0 , 0 TO 0);
		 result : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT or14x16
	PORT(data0x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data10x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data11x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data12x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data13x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data14x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data15x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data4x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data5x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data6x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data7x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data8x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data9x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT reg16nc
	PORT(clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT and14b
	PORT(data0x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	b :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	bb :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	data :  STD_LOGIC_VECTOR(223 DOWNTO 0);
SIGNAL	o :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	or :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	p :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;

SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_2 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_3 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_4 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_5 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_8 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_9 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_10 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_11 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_12 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_13 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_6 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);
SIGNAL	GDFX_TEMP_SIGNAL_7 :  STD_LOGIC_VECTOR(14 DOWNTO 0 , 0 TO 0);

BEGIN 

GDFX_TEMP_SIGNAL_0 <= (b(15 DOWNTO 2) & b(0));
GDFX_TEMP_SIGNAL_1 <= (b(15 DOWNTO 3) & b(1 DOWNTO 0));
GDFX_TEMP_SIGNAL_2 <= (b(15 DOWNTO 4) & b(2 DOWNTO 0));
GDFX_TEMP_SIGNAL_3 <= (b(15 DOWNTO 5) & b(3 DOWNTO 0));
GDFX_TEMP_SIGNAL_4 <= (b(15 DOWNTO 6) & b(4 DOWNTO 0));
GDFX_TEMP_SIGNAL_5 <= (b(15 DOWNTO 7) & b(5 DOWNTO 0));
GDFX_TEMP_SIGNAL_8 <= (b(15 DOWNTO 10) & b(8 DOWNTO 0));
GDFX_TEMP_SIGNAL_9 <= (b(15 DOWNTO 11) & b(9 DOWNTO 0));
GDFX_TEMP_SIGNAL_10 <= (b(15 DOWNTO 12) & b(10 DOWNTO 0));
GDFX_TEMP_SIGNAL_11 <= (b(15 DOWNTO 13) & b(11 DOWNTO 0));
GDFX_TEMP_SIGNAL_12 <= (b(15 DOWNTO 14) & b(12 DOWNTO 0));
GDFX_TEMP_SIGNAL_13 <= (b(15) & b(13 DOWNTO 0));
GDFX_TEMP_SIGNAL_6 <= (b(15 DOWNTO 8) & b(6 DOWNTO 0));
GDFX_TEMP_SIGNAL_7 <= (b(15 DOWNTO 9) & b(7 DOWNTO 0));


b2v_inst : and16
PORT MAP(data0x => SYNTHESIZED_WIRE_94,
		 data1x => compr_mask,
		 result => b);


b2v_inst1 : or16b
PORT MAP(data => or,
		 result => SYNTHESIZED_WIRE_42);


p(4) <= b(4) AND SYNTHESIZED_WIRE_95;


p(5) <= b(5) AND SYNTHESIZED_WIRE_95 AND bb(4);


p(7) <= b(7) AND SYNTHESIZED_WIRE_95 AND SYNTHESIZED_WIRE_4;


b2v_inst13 : and4b
PORT MAP(data => bb(3 DOWNTO 0),
		 result => SYNTHESIZED_WIRE_95);


b2v_inst14 : and3b
PORT MAP(data => bb(2 DOWNTO 0),
		 result => SYNTHESIZED_WIRE_93);


b2v_inst15 : and2b
PORT MAP(data => bb(1 DOWNTO 0),
		 result => SYNTHESIZED_WIRE_84);


p(6) <= b(6) AND SYNTHESIZED_WIRE_95 AND SYNTHESIZED_WIRE_6;


b2v_inst163 : or15b
PORT MAP(data => b(15 DOWNTO 1),
		 result => SYNTHESIZED_WIRE_13);


b2v_inst164 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_0,
		 result => SYNTHESIZED_WIRE_27);


b2v_inst166 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_1,
		 result => SYNTHESIZED_WIRE_15);


b2v_inst168 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_2,
		 result => SYNTHESIZED_WIRE_17);


b2v_inst17 : inv16b
PORT MAP(data => b,
		 result => bb);


b2v_inst170 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_3,
		 result => SYNTHESIZED_WIRE_19);


b2v_inst172 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_4,
		 result => SYNTHESIZED_WIRE_23);


b2v_inst174 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_5,
		 result => SYNTHESIZED_WIRE_25);


b2v_inst176 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_6,
		 result => SYNTHESIZED_WIRE_21);


b2v_inst178 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_7,
		 result => SYNTHESIZED_WIRE_41);


p(8) <= b(8) AND SYNTHESIZED_WIRE_95 AND SYNTHESIZED_WIRE_8;


b2v_inst180 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_8,
		 result => SYNTHESIZED_WIRE_31);


b2v_inst182 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_9,
		 result => SYNTHESIZED_WIRE_29);


b2v_inst184 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_10,
		 result => SYNTHESIZED_WIRE_35);


b2v_inst186 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_11,
		 result => SYNTHESIZED_WIRE_33);


b2v_inst188 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_12,
		 result => SYNTHESIZED_WIRE_39);


p(9) <= b(9) AND SYNTHESIZED_WIRE_96 AND bb(8);


b2v_inst190 : or15b
PORT MAP(data => GDFX_TEMP_SIGNAL_13,
		 result => SYNTHESIZED_WIRE_37);


b2v_inst192 : or15b
PORT MAP(data => b(14 DOWNTO 0),
		 result => SYNTHESIZED_WIRE_46);


b2v_inst199 : inv1
PORT MAP(data => b(1),
		 result => SYNTHESIZED_WIRE_26);

SYNTHESIZED_WIRE_78 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(13);



p(10) <= b(10) AND SYNTHESIZED_WIRE_96 AND SYNTHESIZED_WIRE_11;


b2v_inst200 : inv1
PORT MAP(data => b(0),
		 result => SYNTHESIZED_WIRE_12);


b2v_inst201 : inv1
PORT MAP(data => b(2),
		 result => SYNTHESIZED_WIRE_14);


b2v_inst202 : inv1
PORT MAP(data => b(3),
		 result => SYNTHESIZED_WIRE_16);


or(0) <= NOT(SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13);


b2v_inst204 : inv1
PORT MAP(data => b(6),
		 result => SYNTHESIZED_WIRE_24);


b2v_inst205 : inv1
PORT MAP(data => b(7),
		 result => SYNTHESIZED_WIRE_20);


b2v_inst206 : inv1
PORT MAP(data => b(4),
		 result => SYNTHESIZED_WIRE_18);


b2v_inst207 : inv1
PORT MAP(data => b(5),
		 result => SYNTHESIZED_WIRE_22);


b2v_inst208 : inv1
PORT MAP(data => b(8),
		 result => SYNTHESIZED_WIRE_40);


b2v_inst209 : inv1
PORT MAP(data => b(9),
		 result => SYNTHESIZED_WIRE_30);

SYNTHESIZED_WIRE_87 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(5);



b2v_inst210 : inv1
PORT MAP(data => b(13),
		 result => SYNTHESIZED_WIRE_38);


b2v_inst211 : inv1
PORT MAP(data => b(14),
		 result => SYNTHESIZED_WIRE_36);


b2v_inst212 : inv1
PORT MAP(data => b(15),
		 result => SYNTHESIZED_WIRE_45);


b2v_inst213 : inv1
PORT MAP(data => b(12),
		 result => SYNTHESIZED_WIRE_32);


b2v_inst214 : inv1
PORT MAP(data => b(10),
		 result => SYNTHESIZED_WIRE_28);


b2v_inst215 : inv1
PORT MAP(data => b(11),
		 result => SYNTHESIZED_WIRE_34);


or(2) <= NOT(SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_15);


or(3) <= NOT(SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_17);


or(4) <= NOT(SYNTHESIZED_WIRE_18 OR SYNTHESIZED_WIRE_19);


or(7) <= NOT(SYNTHESIZED_WIRE_20 OR SYNTHESIZED_WIRE_21);


b2v_inst22 : inv16b
PORT MAP(data => p,
		 result => SYNTHESIZED_WIRE_50);


or(5) <= NOT(SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23);


or(6) <= NOT(SYNTHESIZED_WIRE_24 OR SYNTHESIZED_WIRE_25);


or(1) <= NOT(SYNTHESIZED_WIRE_26 OR SYNTHESIZED_WIRE_27);


or(10) <= NOT(SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29);


or(9) <= NOT(SYNTHESIZED_WIRE_30 OR SYNTHESIZED_WIRE_31);


or(12) <= NOT(SYNTHESIZED_WIRE_32 OR SYNTHESIZED_WIRE_33);


or(11) <= NOT(SYNTHESIZED_WIRE_34 OR SYNTHESIZED_WIRE_35);


or(14) <= NOT(SYNTHESIZED_WIRE_36 OR SYNTHESIZED_WIRE_37);


or(13) <= NOT(SYNTHESIZED_WIRE_38 OR SYNTHESIZED_WIRE_39);


or(8) <= NOT(SYNTHESIZED_WIRE_40 OR SYNTHESIZED_WIRE_41);


b2v_inst23 : reg13set
PORT MAP(sset => SYNTHESIZED_WIRE_42,
		 clock => clk,
		 enable => enable,
		 aset => SYNTHESIZED_WIRE_43,
		 data => SYNTHESIZED_WIRE_44,
		 q => SYNTHESIZED_WIRE_94);


or(15) <= NOT(SYNTHESIZED_WIRE_45 OR SYNTHESIZED_WIRE_46);


b2v_inst231 : inv1
PORT MAP(data => reset,
		 result => SYNTHESIZED_WIRE_43);


b2v_inst232 : inv1
PORT MAP(data => SYNTHESIZED_WIRE_47,
		 result => SYNTHESIZED_WIRE_96);


b2v_inst233 : inv1
PORT MAP(data => SYNTHESIZED_WIRE_48,
		 result => SYNTHESIZED_WIRE_97);


b2v_inst24 : and16
PORT MAP(data0x => SYNTHESIZED_WIRE_94,
		 data1x => SYNTHESIZED_WIRE_50,
		 result => SYNTHESIZED_WIRE_44);


p(11) <= b(11) AND SYNTHESIZED_WIRE_96 AND SYNTHESIZED_WIRE_52;


p(12) <= b(12) AND SYNTHESIZED_WIRE_96 AND SYNTHESIZED_WIRE_54;


p(13) <= b(13) AND SYNTHESIZED_WIRE_97 AND bb(12);

SYNTHESIZED_WIRE_79 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(12);


SYNTHESIZED_WIRE_76 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(15);



p(0) <= b(0) AND b(0);

SYNTHESIZED_WIRE_77 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(14);


SYNTHESIZED_WIRE_83 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(8);


SYNTHESIZED_WIRE_80 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(11);


SYNTHESIZED_WIRE_81 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(10);


SYNTHESIZED_WIRE_88 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(4);



b2v_inst35 : and4b
PORT MAP(data => bb(7 DOWNTO 4),
		 result => SYNTHESIZED_WIRE_8);


b2v_inst36 : and3b
PORT MAP(data => bb(6 DOWNTO 4),
		 result => SYNTHESIZED_WIRE_4);


b2v_inst37 : and2b
PORT MAP(data => bb(5 DOWNTO 4),
		 result => SYNTHESIZED_WIRE_6);


b2v_inst38 : and4b
PORT MAP(data => bb(11 DOWNTO 8),
		 result => SYNTHESIZED_WIRE_54);


b2v_inst39 : and3b
PORT MAP(data => bb(10 DOWNTO 8),
		 result => SYNTHESIZED_WIRE_52);


b2v_inst4 : const2
PORT MAP(		 result => o(15 DOWNTO 14));


b2v_inst40 : and2b
PORT MAP(data => bb(9 DOWNTO 8),
		 result => SYNTHESIZED_WIRE_11);


p(14) <= b(14) AND SYNTHESIZED_WIRE_97 AND SYNTHESIZED_WIRE_57;


p(15) <= b(15) AND SYNTHESIZED_WIRE_97 AND SYNTHESIZED_WIRE_59;

SYNTHESIZED_WIRE_85 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(7);



b2v_inst45 : or8b
PORT MAP(data => b(7 DOWNTO 0),
		 result => SYNTHESIZED_WIRE_47);


b2v_inst46 : or12b
PORT MAP(data => b(11 DOWNTO 0),
		 result => SYNTHESIZED_WIRE_48);

SYNTHESIZED_WIRE_86 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(6);


SYNTHESIZED_WIRE_91 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(1);


SYNTHESIZED_WIRE_92 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(0);


SYNTHESIZED_WIRE_82 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(9);


SYNTHESIZED_WIRE_89 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(3);


SYNTHESIZED_WIRE_90 <= (p & p & p & p & p & p & p & p & p & p & p & p & p & p)(2);



b2v_inst55 : and3b
PORT MAP(data => bb(14 DOWNTO 12),
		 result => SYNTHESIZED_WIRE_59);


b2v_inst56 : and2b
PORT MAP(data => bb(13 DOWNTO 12),
		 result => SYNTHESIZED_WIRE_57);


b2v_inst57 : or14x16
PORT MAP(data0x => SYNTHESIZED_WIRE_60,
		 data10x => SYNTHESIZED_WIRE_61,
		 data11x => SYNTHESIZED_WIRE_62,
		 data12x => SYNTHESIZED_WIRE_63,
		 data13x => SYNTHESIZED_WIRE_64,
		 data14x => SYNTHESIZED_WIRE_65,
		 data15x => SYNTHESIZED_WIRE_66,
		 data1x => SYNTHESIZED_WIRE_67,
		 data2x => SYNTHESIZED_WIRE_68,
		 data3x => SYNTHESIZED_WIRE_69,
		 data4x => SYNTHESIZED_WIRE_70,
		 data5x => SYNTHESIZED_WIRE_71,
		 data6x => SYNTHESIZED_WIRE_72,
		 data7x => SYNTHESIZED_WIRE_73,
		 data8x => SYNTHESIZED_WIRE_74,
		 data9x => SYNTHESIZED_WIRE_75,
		 result => o(13 DOWNTO 0));


b2v_inst6 : reg16nc
PORT MAP(clock => clk,
		 data => o,
		 q => out);


p(1) <= b(1) AND bb(0);


b2v_inst72 : and14b
PORT MAP(data0x => data(223 DOWNTO 210),
		 data1x => SYNTHESIZED_WIRE_76,
		 result => SYNTHESIZED_WIRE_60);


b2v_inst73 : and14b
PORT MAP(data0x => data(209 DOWNTO 196),
		 data1x => SYNTHESIZED_WIRE_77,
		 result => SYNTHESIZED_WIRE_67);


b2v_inst74 : and14b
PORT MAP(data0x => data(195 DOWNTO 182),
		 data1x => SYNTHESIZED_WIRE_78,
		 result => SYNTHESIZED_WIRE_68);


b2v_inst75 : and14b
PORT MAP(data0x => data(181 DOWNTO 168),
		 data1x => SYNTHESIZED_WIRE_79,
		 result => SYNTHESIZED_WIRE_69);


b2v_inst76 : and14b
PORT MAP(data0x => data(167 DOWNTO 154),
		 data1x => SYNTHESIZED_WIRE_80,
		 result => SYNTHESIZED_WIRE_70);


b2v_inst77 : and14b
PORT MAP(data0x => data(153 DOWNTO 140),
		 data1x => SYNTHESIZED_WIRE_81,
		 result => SYNTHESIZED_WIRE_71);


b2v_inst78 : and14b
PORT MAP(data0x => data(139 DOWNTO 126),
		 data1x => SYNTHESIZED_WIRE_82,
		 result => SYNTHESIZED_WIRE_72);


b2v_inst79 : and14b
PORT MAP(data0x => data(125 DOWNTO 112),
		 data1x => SYNTHESIZED_WIRE_83,
		 result => SYNTHESIZED_WIRE_73);


p(2) <= b(2) AND SYNTHESIZED_WIRE_84;


b2v_inst80 : and14b
PORT MAP(data0x => data(111 DOWNTO 98),
		 data1x => SYNTHESIZED_WIRE_85,
		 result => SYNTHESIZED_WIRE_74);


b2v_inst81 : and14b
PORT MAP(data0x => data(97 DOWNTO 84),
		 data1x => SYNTHESIZED_WIRE_86,
		 result => SYNTHESIZED_WIRE_75);


b2v_inst82 : and14b
PORT MAP(data0x => data(83 DOWNTO 70),
		 data1x => SYNTHESIZED_WIRE_87,
		 result => SYNTHESIZED_WIRE_61);


b2v_inst83 : and14b
PORT MAP(data0x => data(69 DOWNTO 56),
		 data1x => SYNTHESIZED_WIRE_88,
		 result => SYNTHESIZED_WIRE_62);


b2v_inst84 : and14b
PORT MAP(data0x => data(55 DOWNTO 42),
		 data1x => SYNTHESIZED_WIRE_89,
		 result => SYNTHESIZED_WIRE_63);


b2v_inst85 : and14b
PORT MAP(data0x => data(41 DOWNTO 28),
		 data1x => SYNTHESIZED_WIRE_90,
		 result => SYNTHESIZED_WIRE_64);


b2v_inst86 : and14b
PORT MAP(data0x => data(27 DOWNTO 14),
		 data1x => SYNTHESIZED_WIRE_91,
		 result => SYNTHESIZED_WIRE_65);


b2v_inst87 : and14b
PORT MAP(data0x => data(13 DOWNTO 0),
		 data1x => SYNTHESIZED_WIRE_92,
		 result => SYNTHESIZED_WIRE_66);


p(3) <= b(3) AND SYNTHESIZED_WIRE_93;

data <= buffer_data;

END bdf_type;