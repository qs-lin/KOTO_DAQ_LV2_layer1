-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 9.1 Build 222 10/21/2009 SJ Full Version"
-- CREATED		"Wed Sep 16 11:43:14 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY min_range IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		enable :  IN  STD_LOGIC;
		reset :  IN  STD_LOGIC;
		use_lossless :  IN  STD_LOGIC;
		data :  IN  STD_LOGIC_VECTOR(13 DOWNTO 0);
		min :  OUT  STD_LOGIC_VECTOR(13 DOWNTO 0);
		range :  OUT  STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END min_range;

ARCHITECTURE bdf_type OF min_range IS 

COMPONENT compare14
	PORT(dataa : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 agb : OUT STD_LOGIC;
		 aleb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT ff3
	PORT(data : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 q : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT reg14nc
	PORT(clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const_loss0
	PORT(		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const_loss1
	PORT(		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const_loss3
	PORT(		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const_loss2
	PORT(		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const_loss4
	PORT(		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const_loss5
	PORT(		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const_loss6
	PORT(		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const_loss7
	PORT(		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT reg14en
	PORT(sclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const_loss14
	PORT(		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT and14b
	PORT(data0x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT reg14en_load
	PORT(sset : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT sub14
	PORT(dataa : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	range_ALTERA_SYNTHESIZED[0] :  STD_LOGIC;
SIGNAL	range_ALTERA_SYNTHESIZED[13] :  STD_LOGIC;
SIGNAL	range_ALTERA_SYNTHESIZED[1] :  STD_LOGIC;
SIGNAL	range_ALTERA_SYNTHESIZED[2] :  STD_LOGIC;
SIGNAL	range_ALTERA_SYNTHESIZED[3] :  STD_LOGIC;
SIGNAL	range_ALTERA_SYNTHESIZED[4] :  STD_LOGIC;
SIGNAL	range_ALTERA_SYNTHESIZED[5] :  STD_LOGIC;
SIGNAL	range_ALTERA_SYNTHESIZED[6] :  STD_LOGIC;
SIGNAL	range_ALTERA_SYNTHESIZED[7] :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC_VECTOR(13 DOWNTO 0);


BEGIN 



b2v_inst : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_71,
		 datab => SYNTHESIZED_WIRE_72,
		 agb => SYNTHESIZED_WIRE_16);


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_2 OR reset;


b2v_inst10 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_73,
		 datab => SYNTHESIZED_WIRE_4,
		 agb => SYNTHESIZED_WIRE_63,
		 aleb => SYNTHESIZED_WIRE_62);


b2v_inst11 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_73,
		 datab => SYNTHESIZED_WIRE_6,
		 aleb => SYNTHESIZED_WIRE_64);


b2v_inst12 : ff3
PORT MAP(data => SYNTHESIZED_WIRE_7,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_19);


b2v_inst13 : reg14nc
PORT MAP(clock => clk,
		 data => SYNTHESIZED_WIRE_74,
		 q => SYNTHESIZED_WIRE_32);


b2v_inst14 : ff3
PORT MAP(data => enable,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_75);


b2v_inst15 : const_loss0
PORT MAP(		 result => SYNTHESIZED_WIRE_31);


b2v_inst16 : const_loss1
PORT MAP(		 result => SYNTHESIZED_WIRE_29);


b2v_inst17 : const_loss3
PORT MAP(		 result => SYNTHESIZED_WIRE_25);


b2v_inst18 : const_loss2
PORT MAP(		 result => SYNTHESIZED_WIRE_27);


b2v_inst19 : ff3
PORT MAP(data => SYNTHESIZED_WIRE_9,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_17);


SYNTHESIZED_WIRE_65 <= SYNTHESIZED_WIRE_10 OR reset;


b2v_inst20 : const_loss4
PORT MAP(		 result => SYNTHESIZED_WIRE_23);


b2v_inst21 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_73,
		 datab => SYNTHESIZED_WIRE_12,
		 agb => SYNTHESIZED_WIRE_59,
		 aleb => SYNTHESIZED_WIRE_58);


SYNTHESIZED_WIRE_10 <= SYNTHESIZED_WIRE_75 AND SYNTHESIZED_WIRE_14;


SYNTHESIZED_WIRE_2 <= SYNTHESIZED_WIRE_75 AND SYNTHESIZED_WIRE_16;



b2v_inst25 : ff3
PORT MAP(data => SYNTHESIZED_WIRE_18,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_34);



b2v_inst27 : const_loss5
PORT MAP(		 result => SYNTHESIZED_WIRE_12);


b2v_inst28 : const_loss6
PORT MAP(		 result => SYNTHESIZED_WIRE_70);


b2v_inst29 : const_loss7
PORT MAP(		 result => SYNTHESIZED_WIRE_4);


b2v_inst3 : reg14en
PORT MAP(sclr => reset,
		 clock => clk,
		 enable => SYNTHESIZED_WIRE_20,
		 data => SYNTHESIZED_WIRE_71,
		 q => SYNTHESIZED_WIRE_72);


b2v_inst30 : const_loss14
PORT MAP(		 result => SYNTHESIZED_WIRE_6);


b2v_inst31 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_73,
		 datab => SYNTHESIZED_WIRE_23,
		 agb => SYNTHESIZED_WIRE_57,
		 aleb => SYNTHESIZED_WIRE_56);


b2v_inst32 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_73,
		 datab => SYNTHESIZED_WIRE_25,
		 agb => SYNTHESIZED_WIRE_55,
		 aleb => SYNTHESIZED_WIRE_54);


b2v_inst33 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_73,
		 datab => SYNTHESIZED_WIRE_27,
		 agb => SYNTHESIZED_WIRE_53,
		 aleb => SYNTHESIZED_WIRE_52);


b2v_inst34 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_73,
		 datab => SYNTHESIZED_WIRE_29,
		 agb => SYNTHESIZED_WIRE_51,
		 aleb => SYNTHESIZED_WIRE_50);


b2v_inst35 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_73,
		 datab => SYNTHESIZED_WIRE_31,
		 agb => SYNTHESIZED_WIRE_49,
		 aleb => SYNTHESIZED_WIRE_45);


b2v_inst36 : and14b
PORT MAP(data0x => SYNTHESIZED_WIRE_32,
		 data1x => SYNTHESIZED_WIRE_33,
		 result => min);

SYNTHESIZED_WIRE_33 <= (use_lossless & use_lossless & use_lossless & use_lossless & use_lossless & use_lossless & use_lossless & use_lossless & use_lossless & use_lossless & use_lossless & use_lossless & use_lossless & use_lossless);




b2v_inst39 : ff3
PORT MAP(data => SYNTHESIZED_WIRE_35,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_36);



b2v_inst41 : ff3
PORT MAP(data => SYNTHESIZED_WIRE_37,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_38);



b2v_inst43 : ff3
PORT MAP(data => SYNTHESIZED_WIRE_39,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_40);



b2v_inst45 : ff3
PORT MAP(data => SYNTHESIZED_WIRE_41,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_42);



b2v_inst47 : ff3
PORT MAP(data => SYNTHESIZED_WIRE_43,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_44);



b2v_inst49 : ff3
PORT MAP(data => SYNTHESIZED_WIRE_45,
		 clock => clk,
		 q => SYNTHESIZED_WIRE_48);


b2v_inst5 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_71,
		 datab => SYNTHESIZED_WIRE_74,
		 aleb => SYNTHESIZED_WIRE_14);



SYNTHESIZED_WIRE_43 <= SYNTHESIZED_WIRE_49 AND SYNTHESIZED_WIRE_50;


SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_51 AND SYNTHESIZED_WIRE_52;


SYNTHESIZED_WIRE_39 <= SYNTHESIZED_WIRE_53 AND SYNTHESIZED_WIRE_54;


SYNTHESIZED_WIRE_37 <= SYNTHESIZED_WIRE_55 AND SYNTHESIZED_WIRE_56;


SYNTHESIZED_WIRE_35 <= SYNTHESIZED_WIRE_57 AND SYNTHESIZED_WIRE_58;


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_59 AND SYNTHESIZED_WIRE_60;


SYNTHESIZED_WIRE_7 <= SYNTHESIZED_WIRE_61 AND SYNTHESIZED_WIRE_62;


SYNTHESIZED_WIRE_9 <= SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64;


b2v_inst6 : reg14en_load
PORT MAP(sset => reset,
		 clock => clk,
		 enable => SYNTHESIZED_WIRE_65,
		 data => SYNTHESIZED_WIRE_71,
		 q => SYNTHESIZED_WIRE_74);


b2v_inst7 : sub14
PORT MAP(dataa => SYNTHESIZED_WIRE_72,
		 datab => SYNTHESIZED_WIRE_74,
		 result => SYNTHESIZED_WIRE_73);


b2v_inst8 : reg14nc
PORT MAP(clock => clk,
		 data => data,
		 q => SYNTHESIZED_WIRE_71);


b2v_inst9 : compare14
PORT MAP(dataa => SYNTHESIZED_WIRE_73,
		 datab => SYNTHESIZED_WIRE_70,
		 agb => SYNTHESIZED_WIRE_61,
		 aleb => SYNTHESIZED_WIRE_60);


END bdf_type;