-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 9.1 Build 222 10/21/2009 SJ Full Version"
-- CREATED		"Wed Sep 16 11:29:57 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY uncompressed_read IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		use_lossless :  IN  STD_LOGIC;
		packet_transfer :  IN  STD_LOGIC;
		data_transfer :  IN  STD_LOGIC;
		in :  IN  STD_LOGIC_VECTOR(223 DOWNTO 0);
		out :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END uncompressed_read;

ARCHITECTURE bdf_type OF uncompressed_read IS 

COMPONENT reg112
	PORT(clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(111 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(111 DOWNTO 0)
	);
END COMPONENT;

COMPONENT const2
	PORT(		 result : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT reg16nc
	PORT(clock : IN STD_LOGIC;
		 data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT counter4
	PORT(clock : IN STD_LOGIC;
		 cnt_en : IN STD_LOGIC;
		 aclr : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux224
	PORT(sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(223 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(223 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(223 DOWNTO 0)
	);
END COMPONENT;

COMPONENT decoder_enable
	PORT(data : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 eq0 : OUT STD_LOGIC;
		 eq1 : OUT STD_LOGIC;
		 eq2 : OUT STD_LOGIC;
		 eq3 : OUT STD_LOGIC;
		 eq4 : OUT STD_LOGIC;
		 eq5 : OUT STD_LOGIC;
		 eq6 : OUT STD_LOGIC;
		 eq7 : OUT STD_LOGIC;
		 eq8 : OUT STD_LOGIC;
		 eq9 : OUT STD_LOGIC;
		 eq10 : OUT STD_LOGIC;
		 eq11 : OUT STD_LOGIC;
		 eq12 : OUT STD_LOGIC;
		 eq13 : OUT STD_LOGIC;
		 eq14 : OUT STD_LOGIC;
		 eq15 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT or14x16
	PORT(data0x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data10x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data11x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data12x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data13x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data14x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data15x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data4x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data5x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data6x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data7x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data8x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data9x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

COMPONENT and14b
	PORT(data0x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	cnt :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	d :  STD_LOGIC_VECTOR(223 DOWNTO 0);
SIGNAL	data :  STD_LOGIC_VECTOR(223 DOWNTO 0);
SIGNAL	o :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(111 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(111 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(111 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(111 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC_VECTOR(111 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC_VECTOR(111 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC_VECTOR(111 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC_VECTOR(111 DOWNTO 0);


BEGIN 



b2v_inst : reg112
PORT MAP(clock => clk,
		 data => in(111 DOWNTO 0),
		 q => SYNTHESIZED_WIRE_3);


b2v_inst1 : reg112
PORT MAP(clock => clk,
		 data => in(223 DOWNTO 112),
		 q => SYNTHESIZED_WIRE_37);

SYNTHESIZED_WIRE_41 <= (SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_0);


SYNTHESIZED_WIRE_45 <= (SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_1);



b2v_inst12 : const2
PORT MAP(		 result => o(15 DOWNTO 14));


b2v_inst13 : reg16nc
PORT MAP(clock => clk,
		 data => o,
		 q => out);


SYNTHESIZED_WIRE_2 <= NOT(packet_transfer);



b2v_inst15 : counter4
PORT MAP(clock => clk,
		 cnt_en => data_transfer,
		 aclr => SYNTHESIZED_WIRE_2,
		 q => cnt);


b2v_inst16 : mux224
PORT MAP(sel => use_lossless,
		 data0x => in,
		 data1x => d,
		 result => data);


b2v_inst17 : decoder_enable
PORT MAP(data => cnt(3 DOWNTO 0),
		 eq0 => SYNTHESIZED_WIRE_17,
		 eq1 => SYNTHESIZED_WIRE_16,
		 eq2 => SYNTHESIZED_WIRE_20,
		 eq3 => SYNTHESIZED_WIRE_19,
		 eq4 => SYNTHESIZED_WIRE_12,
		 eq5 => SYNTHESIZED_WIRE_4,
		 eq6 => SYNTHESIZED_WIRE_15,
		 eq7 => SYNTHESIZED_WIRE_14,
		 eq8 => SYNTHESIZED_WIRE_9,
		 eq9 => SYNTHESIZED_WIRE_1,
		 eq10 => SYNTHESIZED_WIRE_11,
		 eq11 => SYNTHESIZED_WIRE_10,
		 eq12 => SYNTHESIZED_WIRE_5,
		 eq13 => SYNTHESIZED_WIRE_0,
		 eq14 => SYNTHESIZED_WIRE_8,
		 eq15 => SYNTHESIZED_WIRE_6);


b2v_inst2 : reg112
PORT MAP(clock => clk,
		 data => SYNTHESIZED_WIRE_3,
		 q => SYNTHESIZED_WIRE_7);

SYNTHESIZED_WIRE_50 <= (SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_4);


SYNTHESIZED_WIRE_42 <= (SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_5);


SYNTHESIZED_WIRE_39 <= (SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_6);



b2v_inst3 : reg112
PORT MAP(clock => clk,
		 data => SYNTHESIZED_WIRE_7,
		 q => SYNTHESIZED_WIRE_13);

SYNTHESIZED_WIRE_40 <= (SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_8);


SYNTHESIZED_WIRE_46 <= (SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_9);


SYNTHESIZED_WIRE_43 <= (SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10 & SYNTHESIZED_WIRE_10);


SYNTHESIZED_WIRE_44 <= (SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_11);


SYNTHESIZED_WIRE_51 <= (SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_12);



b2v_inst4 : reg112
PORT MAP(clock => clk,
		 data => SYNTHESIZED_WIRE_13,
		 q => SYNTHESIZED_WIRE_18);

SYNTHESIZED_WIRE_48 <= (SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14 & SYNTHESIZED_WIRE_14);


SYNTHESIZED_WIRE_49 <= (SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_15);


SYNTHESIZED_WIRE_54 <= (SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_16);


SYNTHESIZED_WIRE_55 <= (SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17);



b2v_inst5 : reg112
PORT MAP(clock => clk,
		 data => SYNTHESIZED_WIRE_18,
		 q => d(111 DOWNTO 0));

SYNTHESIZED_WIRE_52 <= (SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_19);


SYNTHESIZED_WIRE_53 <= (SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_20);



b2v_inst57 : or14x16
PORT MAP(data0x => SYNTHESIZED_WIRE_21,
		 data10x => SYNTHESIZED_WIRE_22,
		 data11x => SYNTHESIZED_WIRE_23,
		 data12x => SYNTHESIZED_WIRE_24,
		 data13x => SYNTHESIZED_WIRE_25,
		 data14x => SYNTHESIZED_WIRE_26,
		 data15x => SYNTHESIZED_WIRE_27,
		 data1x => SYNTHESIZED_WIRE_28,
		 data2x => SYNTHESIZED_WIRE_29,
		 data3x => SYNTHESIZED_WIRE_30,
		 data4x => SYNTHESIZED_WIRE_31,
		 data5x => SYNTHESIZED_WIRE_32,
		 data6x => SYNTHESIZED_WIRE_33,
		 data7x => SYNTHESIZED_WIRE_34,
		 data8x => SYNTHESIZED_WIRE_35,
		 data9x => SYNTHESIZED_WIRE_36,
		 result => o(13 DOWNTO 0));


b2v_inst6 : reg112
PORT MAP(clock => clk,
		 data => SYNTHESIZED_WIRE_37,
		 q => SYNTHESIZED_WIRE_38);


b2v_inst7 : reg112
PORT MAP(clock => clk,
		 data => SYNTHESIZED_WIRE_38,
		 q => SYNTHESIZED_WIRE_47);


b2v_inst72 : and14b
PORT MAP(data0x => data(223 DOWNTO 210),
		 data1x => SYNTHESIZED_WIRE_39,
		 result => SYNTHESIZED_WIRE_21);


b2v_inst73 : and14b
PORT MAP(data0x => data(209 DOWNTO 196),
		 data1x => SYNTHESIZED_WIRE_40,
		 result => SYNTHESIZED_WIRE_28);


b2v_inst74 : and14b
PORT MAP(data0x => data(195 DOWNTO 182),
		 data1x => SYNTHESIZED_WIRE_41,
		 result => SYNTHESIZED_WIRE_29);


b2v_inst75 : and14b
PORT MAP(data0x => data(181 DOWNTO 168),
		 data1x => SYNTHESIZED_WIRE_42,
		 result => SYNTHESIZED_WIRE_30);


b2v_inst76 : and14b
PORT MAP(data0x => data(167 DOWNTO 154),
		 data1x => SYNTHESIZED_WIRE_43,
		 result => SYNTHESIZED_WIRE_31);


b2v_inst77 : and14b
PORT MAP(data0x => data(153 DOWNTO 140),
		 data1x => SYNTHESIZED_WIRE_44,
		 result => SYNTHESIZED_WIRE_32);


b2v_inst78 : and14b
PORT MAP(data0x => data(139 DOWNTO 126),
		 data1x => SYNTHESIZED_WIRE_45,
		 result => SYNTHESIZED_WIRE_33);


b2v_inst79 : and14b
PORT MAP(data0x => data(125 DOWNTO 112),
		 data1x => SYNTHESIZED_WIRE_46,
		 result => SYNTHESIZED_WIRE_34);


b2v_inst8 : reg112
PORT MAP(clock => clk,
		 data => SYNTHESIZED_WIRE_47,
		 q => SYNTHESIZED_WIRE_56);


b2v_inst80 : and14b
PORT MAP(data0x => data(111 DOWNTO 98),
		 data1x => SYNTHESIZED_WIRE_48,
		 result => SYNTHESIZED_WIRE_35);


b2v_inst81 : and14b
PORT MAP(data0x => data(97 DOWNTO 84),
		 data1x => SYNTHESIZED_WIRE_49,
		 result => SYNTHESIZED_WIRE_36);


b2v_inst82 : and14b
PORT MAP(data0x => data(83 DOWNTO 70),
		 data1x => SYNTHESIZED_WIRE_50,
		 result => SYNTHESIZED_WIRE_22);


b2v_inst83 : and14b
PORT MAP(data0x => data(69 DOWNTO 56),
		 data1x => SYNTHESIZED_WIRE_51,
		 result => SYNTHESIZED_WIRE_23);


b2v_inst84 : and14b
PORT MAP(data0x => data(55 DOWNTO 42),
		 data1x => SYNTHESIZED_WIRE_52,
		 result => SYNTHESIZED_WIRE_24);


b2v_inst85 : and14b
PORT MAP(data0x => data(41 DOWNTO 28),
		 data1x => SYNTHESIZED_WIRE_53,
		 result => SYNTHESIZED_WIRE_25);


b2v_inst86 : and14b
PORT MAP(data0x => data(27 DOWNTO 14),
		 data1x => SYNTHESIZED_WIRE_54,
		 result => SYNTHESIZED_WIRE_26);


b2v_inst87 : and14b
PORT MAP(data0x => data(13 DOWNTO 0),
		 data1x => SYNTHESIZED_WIRE_55,
		 result => SYNTHESIZED_WIRE_27);


b2v_inst9 : reg112
PORT MAP(clock => clk,
		 data => SYNTHESIZED_WIRE_56,
		 q => d(223 DOWNTO 112));


END bdf_type;